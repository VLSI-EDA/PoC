-- EMACS settings: -*-  tab-width: 4; indent-tabs-mode: t -*-
-- vim: tabstop=4:shiftwidth=4:noexpandtab
-- kate: tab-width 4; replace-tabs off; indent-width 4;
-- =============================================================================
-- Authors:					Paul Genssler
--
-- Entity:					ICAP Dini PCIe Controller
--
-- Description:
-- -------------------------------------
-- This module was designed to connect the Xilinx "Internal Configuration Access Port" (ICAP)
-- to a PCIe endpoint on a Dini board. Tested on:
--
-- tbd
--
-- License:
-- =============================================================================
-- Copyright 2007-2016 Technische Universitaet Dresden - Germany,
--										 Chair for VLSI-Design, Diagnostics and Architecture
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--		http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
-- =============================================================================
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

library UNISIM;
use UNISIM.vcomponents.all;

library poc;
use poc.utils.all;


entity icap_dini is
	generic (
		CLKIN1_PERIOD	  : real := 8.0;		-- divide input clk
		CLKOUT0_DIVIDE_F  : real := 6.25;		-- multiply to get 100 MHz
		MIN_DEPTH_OUT     : positive := 256;
		MIN_DEPTH_IN      : positive := 256
	);
	port (
		clk 			: in	std_logic;
		res				: in	std_logic;
				
		---- external clock ---- 
		status_in		: in	std_logic_vector(31 downto 0);	
		status_out		: out	std_logic_vector(31 downto 0);
		
		-- data in
		write_put		: in	std_logic;
		write_full		: out	std_logic;
		write_data		: in	std_logic_vector(31 DOWNTO 0);
		
		-- data out
		read_got		: in		std_logic;
		read_full 		: out		std_logic;
		read_data 		: out		std_logic_vector(31 DOWNTO 0)
	);
end icap_dini;

architecture Behavioral of icap_dini is
	signal reset					: std_logic;
	signal icap_clk					: std_logic;
	signal icap_clk_locked			: std_logic;
	signal icap_clk_feedback		: std_logic;
	
	signal status_write_done		: std_logic;
	signal status_write_done_d		: std_logic;
	signal status_write_done_flank	: std_logic;
	signal status_write_done_icapclk: std_logic;

	constant STATUS_PLACES_WRITE_DONE		: natural := 0;
	constant STATUS_PLACES_RESET			: natural := 1;
	constant STATUS_PLACES_PARTIAL_RESET	: natural := 2;
	constant STATUS_PLACES_READBACK			: natural := 3;
	constant STATUS_PLACES_ICAP_ERROR		: natural := 4;
	constant STATUS_PLACES_FSM_IDLE			: natural := 5;

	signal in_data_valid			: std_logic;
	constant STATE_BITS 			: positive := 2;
	constant state_almost_full		: std_logic_vector(STATE_BITS -1 downto 0) := (0 => '0', others => '1');
	signal in_data_fill_state		: std_logic_vector(STATE_BITS -1 downto 0);
	signal in_data_rden				: std_logic;
	signal in_data_start			: std_logic;		-- high after enough data was written into the pci->icap fifo
														--  or write done (status register)
	signal icap_rden				: std_logic;		-- icap wants some yummy data
	signal in_data					: std_logic_vector(31 downto 0);
	
	signal out_data_full			: std_logic;
	signal out_data_put				: std_logic;
	signal out_data					: std_logic_vector(31 downto 0);
	
	signal icap_data_config			: std_logic_vector(31 downto 0);
	signal icap_data_readback		: std_logic_vector(31 downto 0);
	signal icap_csb					: std_logic;
	signal icap_rw					: std_logic;
	
	signal icap_data_config_r		: std_logic_vector(31 downto 0);
	signal icap_data_readback_r		: std_logic_vector(31 downto 0);
	signal icap_csb_r				: std_logic;
	signal icap_rw_r				: std_logic;
	
	signal fsm_status				: std_logic_vector(31 downto 0);
	signal fsm_status_clk			: std_logic_vector(31 downto 0);
	signal fsm_ready				: std_logic;
	signal fsm_ready_d				: std_logic;
begin
	reset <= res or status_in(STATUS_PLACES_RESET) or not icap_clk_locked;
	status_write_done <= status_in(STATUS_PLACES_WRITE_DONE);
	status_write_done_d <= status_write_done when rising_edge(clk);
	status_write_done_flank <= to_sl(status_write_done = '1' and status_write_done_d = '0');
	
	status_out <= (STATUS_PLACES_PARTIAL_RESET	=> fsm_status_clk(0),
					STATUS_PLACES_READBACK		=> fsm_status_clk(1),
					STATUS_PLACES_ICAP_ERROR	=> fsm_status_clk(2),
					STATUS_PLACES_FSM_IDLE		=> fsm_status_clk(3),
					others => '0');
					
	fsm_ready <= fsm_status(3);
	fsm_ready_d <= fsm_ready when rising_edge(icap_clk);

	-- buffer some data before starting the icap, icap needs to be sync'ed before it can be paused
	in_data_buffer_p : process (icap_clk) begin
		if (rising_edge(icap_clk)) then
			if (reset = '1') then
				in_data_start <= '0';
			else
				if fsm_ready = '1' and fsm_ready_d = '0' then	-- reset after icap is done
					in_data_start <= '0';
				elsif in_data_fill_state = state_almost_full or status_write_done_icapclk = '1' then	-- set when fifo almost full or write already done
					in_data_start <= '1';
				end if;
			end if;
		end if;	
	end process in_data_buffer_p;
	
	in_data_rden <= icap_rden and in_data_start and in_data_valid;
		
	-- sync the written pci data into the user clk
	-- writer: pci
	-- reader: core
	fifo_in : ENTITY poc.fifo_ic_got
		generic map(
			D_BITS			=> 32,
			MIN_DEPTH		=> MIN_DEPTH_IN,
			OUTPUT_REG		=> false,
			FSTATE_RD_BITS	=> STATE_BITS
		)
		port map(
			clk_wr 			=> clk,
			rst_wr 			=> reset,
			put    			=> write_put,
			din    			=> write_data,
			full   			=> write_full,
			estate_wr		=> open,

			clk_rd 			=> icap_clk,
			rst_rd 			=> reset,
			got    			=> in_data_rden,
			valid  			=> in_data_valid,
			dout   			=> in_data,
			fstate_rd		=> in_data_fill_state
		);
	
	-- sync data from this core to the pci bus
	-- writer: core
	-- reader: pci
	fifo_out : ENTITY poc.fifo_ic_got
		generic map(
			D_BITS			=> 32,
			MIN_DEPTH		=> MIN_DEPTH_OUT,
			OUTPUT_REG		=> false
		)
		port map(
			clk_wr 			=> icap_clk,
			rst_wr 			=> reset,
			put    			=> out_data_put,
			din    			=> out_data,
			full   			=> out_data_full,

			clk_rd 			=> clk,
			rst_rd 			=> reset,
			got    			=> read_got,
			valid  			=> read_full,
			dout   			=> read_data
		);
		
	icap_fsm_inst: entity work.icap_fsm PORT MAP(
		clk => icap_clk,
		reset => reset,
		icap_in => icap_data_config_r,
		icap_out => icap_data_readback_r,
		icap_csb => icap_csb_r,
		icap_rw => icap_rw_r,
		in_data => in_data,
		in_data_valid => in_data_rden,		-- TODO start one clock cycle later
		in_data_rden => icap_rden,
		out_data => out_data,
		out_data_valid => out_data_put,
		out_data_full => out_data_full,
		status => fsm_status
	);
	
	-- icap
	icap_reg_p : process (icap_clk) begin
		if rising_edge(icap_clk) then
			icap_data_readback_r <= icap_data_readback;
			icap_csb <= icap_csb_r;
			icap_rw <= icap_rw_r;
			icap_data_config <= icap_data_config_r;
		end if;
	end process icap_reg_p;
	
	icap_inst : entity poc.xil_ICAP
	port map (
		clk			=> icap_clk,
		disable		=> icap_csb,
		busy		=> open,
		data_in		=> icap_data_config,
		data_out	=> icap_data_readback,
		rd_wr		=> icap_rw
	);
	
	-- icap clock generation
   MMCME2_BASE_inst : MMCME2_BASE
   generic map (
      BANDWIDTH => "OPTIMIZED",  -- OPTIMIZED, HIGH, LOW
      CLKIN1_PERIOD => CLKIN1_PERIOD,      -- Input clock period in ns to ps resolution (i.e. 33.333 is 30 MHz).
      CLKOUT0_DIVIDE_F => CLKOUT0_DIVIDE_F
   )
   port map (
      -- Clock Outputs: 1-bit (each) output: User configurable clock outputs
      CLKOUT0 => icap_clk,   -- 1-bit output: CLKOUT0
      CLKOUT0B => open,   -- 1-bit output: Inverted CLKOUT0
      CLKOUT1 => open,     -- 1-bit output: CLKOUT1
      CLKOUT1B => open,   -- 1-bit output: Inverted CLKOUT1
      CLKOUT2 => open,     -- 1-bit output: CLKOUT2
      CLKOUT2B => open,   -- 1-bit output: Inverted CLKOUT2
      CLKOUT3 => open,     -- 1-bit output: CLKOUT3
      CLKOUT3B => open,   -- 1-bit output: Inverted CLKOUT3
      CLKOUT4 => open,     -- 1-bit output: CLKOUT4
      CLKOUT5 => open,     -- 1-bit output: CLKOUT5
      CLKOUT6 => open,     -- 1-bit output: CLKOUT6
      -- Feedback Clocks: 1-bit (each) output: Clock feedback ports
      CLKFBOUT => icap_clk_feedback, -- 1-bit output: Feedback clock
      CLKFBOUTB => open,
      LOCKED => icap_clk_locked,     -- 1-bit output: LOCK
      CLKIN1 => clk,     -- 1-bit input: Input clock
      -- Control Ports: 1-bit (each) input: PLL control ports
      PWRDWN => '0',     -- 1-bit input: Power-down
      RST => '0',           -- 1-bit input: Reset
      -- Feedback Clocks: 1-bit (each) input: Clock feedback ports
      CLKFBIN => icap_clk_feedback    -- 1-bit input: Feedback clock
   );
	
	bit_sync : entity poc.sync_Strobe
	port map (
		clock1 => clk,
		clock2 => icap_clk,
		input(0) => status_write_done_flank,
		output(0) => status_write_done_icapclk,
		busy => open
	);
	
	fsm_status_sync : entity poc.sync_vector
	generic map (
		master_bits => 32
	) port map (
		clock1 => icap_clk,
		clock2 => clk,
		input => fsm_status,
		output => fsm_status_clk,
		busy => open,
		changed => open
	);
	
	
end Behavioral;
